`define WIDTH 8

`define NEW_OBJ\
function new(string name="");\
	super.new(name);\
endfunction

`define NEW_COMP\
function new(string name="" ,uvm_component parent);\
	super.new(name,parent);\
endfunction

uvm_factory factory= uvm_factory::get();
