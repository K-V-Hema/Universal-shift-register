typedef uvm_sequencer #(usr_tx)usr_sqr;
